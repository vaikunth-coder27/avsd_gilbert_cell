magic
tech sky130A
timestamp 1629118681
<< nmos >>
rect 45 0 63 600
rect 213 0 231 600
rect 376 0 394 600
rect 544 0 562 600
<< ndiff >>
rect 0 563 45 600
rect 0 546 14 563
rect 32 546 45 563
rect 0 529 45 546
rect 0 512 14 529
rect 32 512 45 529
rect 0 490 45 512
rect 0 473 14 490
rect 32 473 45 490
rect 0 451 45 473
rect 0 434 14 451
rect 32 434 45 451
rect 0 412 45 434
rect 0 395 14 412
rect 32 395 45 412
rect 0 378 45 395
rect 0 361 14 378
rect 32 361 45 378
rect 0 344 45 361
rect 0 327 14 344
rect 32 327 45 344
rect 0 310 45 327
rect 0 293 14 310
rect 32 293 45 310
rect 0 272 45 293
rect 0 255 14 272
rect 32 255 45 272
rect 0 238 45 255
rect 0 221 14 238
rect 32 221 45 238
rect 0 204 45 221
rect 0 187 14 204
rect 32 187 45 204
rect 0 170 45 187
rect 0 153 14 170
rect 32 153 45 170
rect 0 136 45 153
rect 0 119 14 136
rect 32 119 45 136
rect 0 102 45 119
rect 0 85 14 102
rect 32 85 45 102
rect 0 67 45 85
rect 0 50 14 67
rect 32 50 45 67
rect 0 32 45 50
rect 0 15 14 32
rect 32 15 45 32
rect 0 0 45 15
rect 63 563 108 600
rect 63 546 77 563
rect 95 546 108 563
rect 63 529 108 546
rect 63 512 77 529
rect 95 512 108 529
rect 63 490 108 512
rect 63 473 77 490
rect 95 473 108 490
rect 63 451 108 473
rect 63 434 77 451
rect 95 434 108 451
rect 63 412 108 434
rect 63 395 77 412
rect 95 395 108 412
rect 63 378 108 395
rect 63 361 77 378
rect 95 361 108 378
rect 63 344 108 361
rect 63 327 77 344
rect 95 327 108 344
rect 63 310 108 327
rect 63 293 77 310
rect 95 293 108 310
rect 63 272 108 293
rect 63 255 77 272
rect 95 255 108 272
rect 63 238 108 255
rect 63 221 77 238
rect 95 221 108 238
rect 63 204 108 221
rect 63 187 77 204
rect 95 187 108 204
rect 63 170 108 187
rect 63 153 77 170
rect 95 153 108 170
rect 63 136 108 153
rect 63 119 77 136
rect 95 119 108 136
rect 63 102 108 119
rect 63 85 77 102
rect 95 85 108 102
rect 63 67 108 85
rect 63 50 77 67
rect 95 50 108 67
rect 63 32 108 50
rect 63 15 77 32
rect 95 15 108 32
rect 63 0 108 15
rect 168 563 213 600
rect 168 546 184 563
rect 202 546 213 563
rect 168 529 213 546
rect 168 512 184 529
rect 202 512 213 529
rect 168 490 213 512
rect 168 473 184 490
rect 202 473 213 490
rect 168 451 213 473
rect 168 434 184 451
rect 202 434 213 451
rect 168 412 213 434
rect 168 395 184 412
rect 202 395 213 412
rect 168 378 213 395
rect 168 361 184 378
rect 202 361 213 378
rect 168 344 213 361
rect 168 327 184 344
rect 202 327 213 344
rect 168 310 213 327
rect 168 293 184 310
rect 202 293 213 310
rect 168 272 213 293
rect 168 255 184 272
rect 202 255 213 272
rect 168 238 213 255
rect 168 221 184 238
rect 202 221 213 238
rect 168 204 213 221
rect 168 187 184 204
rect 202 187 213 204
rect 168 170 213 187
rect 168 153 184 170
rect 202 153 213 170
rect 168 136 213 153
rect 168 119 184 136
rect 202 119 213 136
rect 168 102 213 119
rect 168 85 184 102
rect 202 85 213 102
rect 168 67 213 85
rect 168 50 184 67
rect 202 50 213 67
rect 168 32 213 50
rect 168 15 184 32
rect 202 15 213 32
rect 168 0 213 15
rect 231 563 276 600
rect 231 546 245 563
rect 263 546 276 563
rect 231 529 276 546
rect 231 512 245 529
rect 263 512 276 529
rect 231 490 276 512
rect 231 473 245 490
rect 263 473 276 490
rect 231 451 276 473
rect 231 434 245 451
rect 263 434 276 451
rect 231 412 276 434
rect 231 395 245 412
rect 263 395 276 412
rect 231 378 276 395
rect 231 361 245 378
rect 263 361 276 378
rect 231 344 276 361
rect 231 327 245 344
rect 263 327 276 344
rect 231 310 276 327
rect 231 293 245 310
rect 263 293 276 310
rect 231 272 276 293
rect 231 255 245 272
rect 263 255 276 272
rect 231 238 276 255
rect 231 221 245 238
rect 263 221 276 238
rect 231 204 276 221
rect 231 187 245 204
rect 263 187 276 204
rect 231 170 276 187
rect 231 153 245 170
rect 263 153 276 170
rect 231 136 276 153
rect 231 119 245 136
rect 263 119 276 136
rect 231 102 276 119
rect 231 85 245 102
rect 263 85 276 102
rect 231 67 276 85
rect 231 50 245 67
rect 263 50 276 67
rect 231 32 276 50
rect 231 15 245 32
rect 263 15 276 32
rect 231 0 276 15
rect 331 563 376 600
rect 331 546 344 563
rect 362 546 376 563
rect 331 529 376 546
rect 331 512 346 529
rect 364 512 376 529
rect 331 490 376 512
rect 331 473 346 490
rect 364 473 376 490
rect 331 451 376 473
rect 331 434 346 451
rect 364 434 376 451
rect 331 412 376 434
rect 331 395 346 412
rect 364 395 376 412
rect 331 378 376 395
rect 331 361 346 378
rect 364 361 376 378
rect 331 344 376 361
rect 331 327 346 344
rect 364 327 376 344
rect 331 310 376 327
rect 331 293 346 310
rect 364 293 376 310
rect 331 272 376 293
rect 331 255 346 272
rect 364 255 376 272
rect 331 238 376 255
rect 331 221 346 238
rect 364 221 376 238
rect 331 204 376 221
rect 331 187 346 204
rect 364 187 376 204
rect 331 170 376 187
rect 331 153 346 170
rect 364 153 376 170
rect 331 136 376 153
rect 331 119 346 136
rect 364 119 376 136
rect 331 102 376 119
rect 331 85 346 102
rect 364 85 376 102
rect 331 67 376 85
rect 331 50 346 67
rect 364 50 376 67
rect 331 32 376 50
rect 331 15 346 32
rect 364 15 376 32
rect 331 0 376 15
rect 394 564 439 600
rect 394 547 408 564
rect 426 547 439 564
rect 394 530 439 547
rect 394 513 408 530
rect 426 513 439 530
rect 394 491 439 513
rect 394 474 408 491
rect 426 474 439 491
rect 394 452 439 474
rect 394 435 408 452
rect 426 435 439 452
rect 394 413 439 435
rect 394 396 408 413
rect 426 396 439 413
rect 394 379 439 396
rect 394 362 408 379
rect 426 362 439 379
rect 394 345 439 362
rect 394 328 408 345
rect 426 328 439 345
rect 394 311 439 328
rect 394 294 408 311
rect 426 294 439 311
rect 394 273 439 294
rect 394 256 408 273
rect 426 256 439 273
rect 394 239 439 256
rect 394 222 408 239
rect 426 222 439 239
rect 394 205 439 222
rect 394 188 408 205
rect 426 188 439 205
rect 394 171 439 188
rect 394 154 408 171
rect 426 154 439 171
rect 394 137 439 154
rect 394 120 408 137
rect 426 120 439 137
rect 394 103 439 120
rect 394 86 408 103
rect 426 86 439 103
rect 394 68 439 86
rect 394 51 408 68
rect 426 51 439 68
rect 394 33 439 51
rect 394 16 408 33
rect 426 16 439 33
rect 394 0 439 16
rect 499 563 544 600
rect 499 546 514 563
rect 532 546 544 563
rect 499 529 544 546
rect 499 512 514 529
rect 532 512 544 529
rect 499 490 544 512
rect 499 473 514 490
rect 532 473 544 490
rect 499 451 544 473
rect 499 434 514 451
rect 532 434 544 451
rect 499 412 544 434
rect 499 395 514 412
rect 532 395 544 412
rect 499 378 544 395
rect 499 361 514 378
rect 532 361 544 378
rect 499 344 544 361
rect 499 327 514 344
rect 532 327 544 344
rect 499 310 544 327
rect 499 293 514 310
rect 532 293 544 310
rect 499 272 544 293
rect 499 255 514 272
rect 532 255 544 272
rect 499 238 544 255
rect 499 221 514 238
rect 532 221 544 238
rect 499 204 544 221
rect 499 187 514 204
rect 532 187 544 204
rect 499 170 544 187
rect 499 153 514 170
rect 532 153 544 170
rect 499 136 544 153
rect 499 119 514 136
rect 532 119 544 136
rect 499 102 544 119
rect 499 85 514 102
rect 532 85 544 102
rect 499 67 544 85
rect 499 50 514 67
rect 532 50 544 67
rect 499 32 544 50
rect 499 15 514 32
rect 532 15 544 32
rect 499 0 544 15
rect 562 564 607 600
rect 562 547 581 564
rect 599 547 607 564
rect 562 530 607 547
rect 562 513 581 530
rect 599 513 607 530
rect 562 491 607 513
rect 562 474 581 491
rect 599 474 607 491
rect 562 452 607 474
rect 562 435 581 452
rect 599 435 607 452
rect 562 413 607 435
rect 562 396 581 413
rect 599 396 607 413
rect 562 379 607 396
rect 562 362 581 379
rect 599 362 607 379
rect 562 345 607 362
rect 562 328 581 345
rect 599 328 607 345
rect 562 311 607 328
rect 562 294 581 311
rect 599 294 607 311
rect 562 273 607 294
rect 562 256 581 273
rect 599 256 607 273
rect 562 239 607 256
rect 562 222 581 239
rect 599 222 607 239
rect 562 205 607 222
rect 562 188 581 205
rect 599 188 607 205
rect 562 171 607 188
rect 562 154 581 171
rect 599 154 607 171
rect 562 137 607 154
rect 562 120 581 137
rect 599 120 607 137
rect 562 103 607 120
rect 562 86 581 103
rect 599 86 607 103
rect 562 68 607 86
rect 562 51 581 68
rect 599 51 607 68
rect 562 33 607 51
rect 562 16 581 33
rect 599 16 607 33
rect 562 0 607 16
<< ndiffc >>
rect 14 797 32 814
rect 578 797 596 814
rect 14 735 32 752
rect 578 735 596 752
rect 14 546 32 563
rect 14 512 32 529
rect 14 473 32 490
rect 14 434 32 451
rect 14 395 32 412
rect 14 361 32 378
rect 14 327 32 344
rect 14 293 32 310
rect 14 255 32 272
rect 14 221 32 238
rect 14 187 32 204
rect 14 153 32 170
rect 14 119 32 136
rect 14 85 32 102
rect 14 50 32 67
rect 14 15 32 32
rect 77 546 95 563
rect 77 512 95 529
rect 77 473 95 490
rect 77 434 95 451
rect 77 395 95 412
rect 77 361 95 378
rect 77 327 95 344
rect 77 293 95 310
rect 77 255 95 272
rect 77 221 95 238
rect 77 187 95 204
rect 77 153 95 170
rect 77 119 95 136
rect 77 85 95 102
rect 77 50 95 67
rect 77 15 95 32
rect 184 546 202 563
rect 184 512 202 529
rect 184 473 202 490
rect 184 434 202 451
rect 184 395 202 412
rect 184 361 202 378
rect 184 327 202 344
rect 184 293 202 310
rect 184 255 202 272
rect 184 221 202 238
rect 184 187 202 204
rect 184 153 202 170
rect 184 119 202 136
rect 184 85 202 102
rect 184 50 202 67
rect 184 15 202 32
rect 245 546 263 563
rect 245 512 263 529
rect 245 473 263 490
rect 245 434 263 451
rect 245 395 263 412
rect 245 361 263 378
rect 245 327 263 344
rect 245 293 263 310
rect 245 255 263 272
rect 245 221 263 238
rect 245 187 263 204
rect 245 153 263 170
rect 245 119 263 136
rect 245 85 263 102
rect 245 50 263 67
rect 245 15 263 32
rect 344 546 362 563
rect 346 512 364 529
rect 346 473 364 490
rect 346 434 364 451
rect 346 395 364 412
rect 346 361 364 378
rect 346 327 364 344
rect 346 293 364 310
rect 346 255 364 272
rect 346 221 364 238
rect 346 187 364 204
rect 346 153 364 170
rect 346 119 364 136
rect 346 85 364 102
rect 346 50 364 67
rect 346 15 364 32
rect 408 547 426 564
rect 408 513 426 530
rect 408 474 426 491
rect 408 435 426 452
rect 408 396 426 413
rect 408 362 426 379
rect 408 328 426 345
rect 408 294 426 311
rect 408 256 426 273
rect 408 222 426 239
rect 408 188 426 205
rect 408 154 426 171
rect 408 120 426 137
rect 408 86 426 103
rect 408 51 426 68
rect 408 16 426 33
rect 514 546 532 563
rect 514 512 532 529
rect 514 473 532 490
rect 514 434 532 451
rect 514 395 532 412
rect 514 361 532 378
rect 514 327 532 344
rect 514 293 532 310
rect 514 255 532 272
rect 514 221 532 238
rect 514 187 532 204
rect 514 153 532 170
rect 514 119 532 136
rect 514 85 532 102
rect 514 50 532 67
rect 514 15 532 32
rect 581 547 599 564
rect 581 513 599 530
rect 581 474 599 491
rect 581 435 599 452
rect 581 396 599 413
rect 581 362 599 379
rect 581 328 599 345
rect 581 294 599 311
rect 581 256 599 273
rect 581 222 599 239
rect 581 188 599 205
rect 581 154 599 171
rect 581 120 599 137
rect 581 86 599 103
rect 581 51 599 68
rect 581 16 599 33
<< psubdiff >>
rect 123 739 166 753
rect 123 722 135 739
rect 154 722 166 739
rect 123 706 166 722
<< psubdiffcont >>
rect 135 722 154 739
<< poly >>
rect 45 600 63 624
rect 213 600 231 624
rect 376 600 394 624
rect 544 600 562 624
rect 45 -15 63 0
rect 213 -15 231 0
rect 376 -15 394 0
rect 544 -15 562 0
rect 37 -20 71 -15
rect 37 -37 45 -20
rect 63 -37 71 -20
rect 37 -45 71 -37
rect 205 -20 239 -15
rect 205 -37 213 -20
rect 231 -37 239 -20
rect 205 -45 239 -37
rect 368 -20 402 -15
rect 368 -37 376 -20
rect 394 -37 402 -20
rect 368 -45 402 -37
rect 536 -20 570 -15
rect 536 -37 544 -20
rect 562 -37 570 -20
rect 536 -45 570 -37
<< polycont >>
rect 45 -37 63 -20
rect 213 -37 231 -20
rect 376 -37 394 -20
rect 544 -37 562 -20
<< ndiffres >>
rect 6 814 39 822
rect 6 797 14 814
rect 32 797 39 814
rect 6 789 39 797
rect 570 814 603 822
rect 570 797 578 814
rect 596 797 603 814
rect 570 789 603 797
rect 14 760 32 789
rect 578 760 596 789
rect 6 752 39 760
rect 6 735 14 752
rect 32 735 39 752
rect 6 727 39 735
rect 570 752 603 760
rect 570 735 578 752
rect 596 735 603 752
rect 570 727 603 735
<< locali >>
rect 6 814 39 822
rect 265 814 322 827
rect 570 814 603 822
rect 6 797 14 814
rect 32 811 578 814
rect 32 797 284 811
rect 6 796 284 797
rect 6 789 39 796
rect 265 794 284 796
rect 302 797 578 811
rect 596 797 603 814
rect 302 796 603 797
rect 302 794 322 796
rect 265 784 322 794
rect 570 789 603 796
rect 6 752 39 760
rect 6 735 14 752
rect 32 735 39 752
rect 6 727 39 735
rect 123 739 166 753
rect 13 589 33 727
rect 123 722 135 739
rect 154 722 166 739
rect 570 752 603 760
rect 570 735 578 752
rect 596 735 603 752
rect 570 727 603 735
rect 123 706 166 722
rect 577 705 597 727
rect 240 679 603 705
rect 240 589 266 679
rect 577 590 603 679
rect 6 569 37 589
rect -57 564 37 569
rect -57 547 -39 564
rect -21 563 37 564
rect -21 547 14 563
rect -57 546 14 547
rect 32 546 37 563
rect -57 541 37 546
rect 6 529 37 541
rect 6 512 14 529
rect 32 512 37 529
rect 6 490 37 512
rect 6 473 14 490
rect 32 473 37 490
rect 6 451 37 473
rect 6 434 14 451
rect 32 434 37 451
rect 6 412 37 434
rect 6 395 14 412
rect 32 395 37 412
rect 6 378 37 395
rect 6 361 14 378
rect 32 361 37 378
rect 6 344 37 361
rect 6 327 14 344
rect 32 327 37 344
rect 6 310 37 327
rect 6 293 14 310
rect 32 293 37 310
rect 6 272 37 293
rect 6 255 14 272
rect 32 255 37 272
rect 6 238 37 255
rect 6 221 14 238
rect 32 221 37 238
rect 6 204 37 221
rect 6 187 14 204
rect 32 187 37 204
rect 6 170 37 187
rect 6 153 14 170
rect 32 153 37 170
rect 6 136 37 153
rect 6 119 14 136
rect 32 119 37 136
rect 6 102 37 119
rect 6 85 14 102
rect 32 85 37 102
rect 6 67 37 85
rect 6 50 14 67
rect 32 50 37 67
rect 6 32 37 50
rect 6 15 14 32
rect 32 15 37 32
rect 6 5 37 15
rect 69 563 100 589
rect 69 546 77 563
rect 95 546 100 563
rect 69 529 100 546
rect 69 512 77 529
rect 95 512 100 529
rect 69 490 100 512
rect 69 473 77 490
rect 95 473 100 490
rect 69 451 100 473
rect 69 434 77 451
rect 95 434 100 451
rect 69 412 100 434
rect 69 395 77 412
rect 95 395 100 412
rect 69 378 100 395
rect 69 361 77 378
rect 95 361 100 378
rect 69 344 100 361
rect 69 327 77 344
rect 95 327 100 344
rect 69 310 100 327
rect 69 293 77 310
rect 95 293 100 310
rect 69 272 100 293
rect 69 255 77 272
rect 95 255 100 272
rect 69 238 100 255
rect 69 221 77 238
rect 95 221 100 238
rect 69 204 100 221
rect 69 187 77 204
rect 95 187 100 204
rect 69 170 100 187
rect 69 153 77 170
rect 95 153 100 170
rect 69 136 100 153
rect 69 119 77 136
rect 95 119 100 136
rect 69 102 100 119
rect 69 85 77 102
rect 95 85 100 102
rect 69 67 100 85
rect 69 50 77 67
rect 95 50 100 67
rect 69 32 100 50
rect 176 563 207 589
rect 238 563 268 589
rect 176 546 184 563
rect 202 546 207 563
rect 176 529 207 546
rect 176 512 184 529
rect 202 512 207 529
rect 176 490 207 512
rect 176 473 184 490
rect 202 473 207 490
rect 176 451 207 473
rect 176 434 184 451
rect 202 434 207 451
rect 176 412 207 434
rect 176 395 184 412
rect 202 395 207 412
rect 176 378 207 395
rect 176 361 184 378
rect 202 361 207 378
rect 176 344 207 361
rect 176 327 184 344
rect 202 327 207 344
rect 176 310 207 327
rect 176 293 184 310
rect 202 293 207 310
rect 176 272 207 293
rect 176 255 184 272
rect 202 255 207 272
rect 176 238 207 255
rect 176 221 184 238
rect 202 221 207 238
rect 176 204 207 221
rect 176 187 184 204
rect 202 187 207 204
rect 176 170 207 187
rect 176 153 184 170
rect 202 153 207 170
rect 176 136 207 153
rect 176 119 184 136
rect 202 119 207 136
rect 176 102 207 119
rect 176 85 184 102
rect 202 85 207 102
rect 176 67 207 85
rect 176 50 184 67
rect 202 50 207 67
rect 176 32 207 50
rect 69 15 77 32
rect 95 15 184 32
rect 202 15 207 32
rect 69 5 100 15
rect 37 -20 71 -15
rect 37 -37 45 -20
rect 63 -37 71 -20
rect 37 -45 71 -37
rect 126 -44 147 15
rect 176 5 207 15
rect 237 546 245 563
rect 263 546 268 563
rect 237 529 268 546
rect 237 512 245 529
rect 263 512 268 529
rect 237 490 268 512
rect 237 473 245 490
rect 263 473 268 490
rect 237 451 268 473
rect 237 434 245 451
rect 263 434 268 451
rect 237 412 268 434
rect 237 395 245 412
rect 263 395 268 412
rect 237 378 268 395
rect 237 361 245 378
rect 263 361 268 378
rect 237 344 268 361
rect 237 327 245 344
rect 263 327 268 344
rect 237 310 268 327
rect 237 293 245 310
rect 263 293 268 310
rect 237 272 268 293
rect 237 255 245 272
rect 263 255 268 272
rect 237 238 268 255
rect 237 221 245 238
rect 263 221 268 238
rect 237 204 268 221
rect 237 187 245 204
rect 263 187 268 204
rect 237 170 268 187
rect 237 153 245 170
rect 263 153 268 170
rect 237 136 268 153
rect 237 119 245 136
rect 263 119 268 136
rect 237 102 268 119
rect 237 85 245 102
rect 263 85 268 102
rect 237 67 268 85
rect 237 50 245 67
rect 263 50 268 67
rect 237 32 268 50
rect 237 15 245 32
rect 263 15 268 32
rect 237 5 268 15
rect 338 563 369 589
rect 338 546 344 563
rect 362 546 369 563
rect 338 529 369 546
rect 338 512 346 529
rect 364 512 369 529
rect 338 490 369 512
rect 338 473 346 490
rect 364 473 369 490
rect 338 451 369 473
rect 338 434 346 451
rect 364 434 369 451
rect 338 412 369 434
rect 338 395 346 412
rect 364 395 369 412
rect 338 378 369 395
rect 338 361 346 378
rect 364 361 369 378
rect 338 344 369 361
rect 338 327 346 344
rect 364 327 369 344
rect 338 310 369 327
rect 338 293 346 310
rect 364 293 369 310
rect 338 272 369 293
rect 338 255 346 272
rect 364 255 369 272
rect 338 238 369 255
rect 338 221 346 238
rect 364 221 369 238
rect 338 204 369 221
rect 338 187 346 204
rect 364 187 369 204
rect 338 170 369 187
rect 338 153 346 170
rect 364 153 369 170
rect 338 136 369 153
rect 338 119 346 136
rect 364 119 369 136
rect 338 102 369 119
rect 338 85 346 102
rect 364 85 369 102
rect 338 67 369 85
rect 338 50 346 67
rect 364 50 369 67
rect 338 32 369 50
rect 338 15 346 32
rect 364 15 369 32
rect 338 5 369 15
rect 400 564 431 590
rect 400 547 408 564
rect 426 547 431 564
rect 400 530 431 547
rect 400 513 408 530
rect 426 513 431 530
rect 400 491 431 513
rect 400 474 408 491
rect 426 474 431 491
rect 400 452 431 474
rect 400 435 408 452
rect 426 435 431 452
rect 400 413 431 435
rect 400 396 408 413
rect 426 396 431 413
rect 400 379 431 396
rect 400 362 408 379
rect 426 362 431 379
rect 400 345 431 362
rect 400 328 408 345
rect 426 328 431 345
rect 400 311 431 328
rect 400 294 408 311
rect 426 294 431 311
rect 400 273 431 294
rect 400 256 408 273
rect 426 256 431 273
rect 400 239 431 256
rect 400 222 408 239
rect 426 222 431 239
rect 400 205 431 222
rect 400 188 408 205
rect 426 188 431 205
rect 400 171 431 188
rect 400 154 408 171
rect 426 154 431 171
rect 400 137 431 154
rect 400 120 408 137
rect 426 120 431 137
rect 400 103 431 120
rect 400 86 408 103
rect 426 86 431 103
rect 400 68 431 86
rect 400 51 408 68
rect 426 51 431 68
rect 400 33 431 51
rect 506 563 537 589
rect 506 546 514 563
rect 532 546 537 563
rect 506 529 537 546
rect 506 512 514 529
rect 532 512 537 529
rect 506 490 537 512
rect 506 473 514 490
rect 532 473 537 490
rect 506 451 537 473
rect 506 434 514 451
rect 532 434 537 451
rect 506 412 537 434
rect 506 395 514 412
rect 532 395 537 412
rect 506 378 537 395
rect 506 361 514 378
rect 532 361 537 378
rect 506 344 537 361
rect 506 327 514 344
rect 532 327 537 344
rect 506 310 537 327
rect 506 293 514 310
rect 532 293 537 310
rect 506 272 537 293
rect 506 255 514 272
rect 532 255 537 272
rect 506 238 537 255
rect 506 221 514 238
rect 532 221 537 238
rect 506 204 537 221
rect 506 187 514 204
rect 532 187 537 204
rect 506 170 537 187
rect 506 153 514 170
rect 532 153 537 170
rect 506 136 537 153
rect 506 119 514 136
rect 532 119 537 136
rect 506 102 537 119
rect 506 85 514 102
rect 532 85 537 102
rect 506 67 537 85
rect 506 50 514 67
rect 532 50 537 67
rect 506 33 537 50
rect 400 16 408 33
rect 426 32 537 33
rect 426 16 514 32
rect 400 6 431 16
rect 205 -19 239 -15
rect 368 -19 402 -15
rect 205 -20 402 -19
rect 205 -37 213 -20
rect 231 -35 376 -20
rect 231 -36 296 -35
rect 231 -37 239 -36
rect 42 -113 65 -45
rect 113 -50 165 -44
rect 205 -45 239 -37
rect 113 -67 130 -50
rect 148 -67 165 -50
rect 113 -84 165 -67
rect 279 -52 296 -36
rect 314 -36 376 -35
rect 314 -52 331 -36
rect 368 -37 376 -36
rect 394 -37 402 -20
rect 368 -45 402 -37
rect 460 -42 481 16
rect 506 15 514 16
rect 532 15 537 32
rect 506 5 537 15
rect 573 569 604 590
rect 573 564 663 569
rect 573 547 581 564
rect 599 547 631 564
rect 649 547 663 564
rect 573 541 663 547
rect 573 530 604 541
rect 573 513 581 530
rect 599 513 604 530
rect 573 491 604 513
rect 573 474 581 491
rect 599 474 604 491
rect 573 452 604 474
rect 573 435 581 452
rect 599 435 604 452
rect 573 413 604 435
rect 573 396 581 413
rect 599 396 604 413
rect 573 379 604 396
rect 573 362 581 379
rect 599 362 604 379
rect 573 345 604 362
rect 573 328 581 345
rect 599 328 604 345
rect 573 311 604 328
rect 573 294 581 311
rect 599 294 604 311
rect 573 273 604 294
rect 573 256 581 273
rect 599 256 604 273
rect 573 239 604 256
rect 573 222 581 239
rect 599 222 604 239
rect 573 205 604 222
rect 573 188 581 205
rect 599 188 604 205
rect 573 171 604 188
rect 573 154 581 171
rect 599 154 604 171
rect 573 137 604 154
rect 573 120 581 137
rect 599 120 604 137
rect 573 103 604 120
rect 573 86 581 103
rect 599 86 604 103
rect 573 68 604 86
rect 573 51 581 68
rect 599 51 604 68
rect 573 33 604 51
rect 573 16 581 33
rect 599 16 604 33
rect 573 6 604 16
rect 536 -20 570 -15
rect 536 -37 544 -20
rect 562 -37 570 -20
rect 279 -70 331 -52
rect 447 -48 498 -42
rect 536 -45 570 -37
rect 447 -65 464 -48
rect 482 -65 498 -48
rect 447 -81 498 -65
rect 543 -113 564 -45
rect 42 -130 564 -113
rect 42 -136 297 -130
rect 279 -137 297 -136
rect 280 -147 297 -137
rect 315 -136 564 -130
rect 315 -137 333 -136
rect 315 -147 332 -137
rect 280 -171 332 -147
<< viali >>
rect 284 794 302 811
rect 135 722 154 739
rect -39 547 -21 564
rect 14 546 32 563
rect 344 546 362 563
rect 130 -67 148 -50
rect 296 -52 314 -35
rect 631 547 649 564
rect 464 -65 482 -48
rect 297 -147 315 -130
<< metal1 >>
rect 265 811 322 827
rect 265 794 284 811
rect 302 794 322 811
rect 265 784 322 794
rect 123 739 166 753
rect 123 722 135 739
rect 154 722 166 739
rect 123 706 166 722
rect 341 569 366 572
rect -57 564 35 569
rect -57 547 -39 564
rect -21 563 35 564
rect 341 563 368 569
rect -21 547 14 563
rect -57 546 14 547
rect 32 546 344 563
rect 362 546 368 563
rect -57 545 368 546
rect -57 541 35 545
rect 341 541 368 545
rect 624 564 663 569
rect 624 547 631 564
rect 649 547 663 564
rect 624 541 663 547
rect 341 540 366 541
rect 286 -35 323 -29
rect 120 -50 157 -44
rect 120 -67 130 -50
rect 148 -67 157 -50
rect 120 -84 157 -67
rect 286 -52 296 -35
rect 314 -52 323 -35
rect 286 -68 323 -52
rect 454 -48 491 -42
rect 454 -65 464 -48
rect 482 -65 491 -48
rect 454 -80 491 -65
rect 287 -130 324 -124
rect 287 -147 297 -130
rect 315 -147 324 -130
rect 287 -167 324 -147
<< labels >>
flabel metal1 136 716 153 719 0 FreeSans 56 0 0 -56 GND
flabel metal1 284 813 302 815 0 FreeSans 56 0 0 56 VDD
flabel metal1 130 -72 148 -70 0 FreeSans 56 0 0 -56 V1
flabel metal1 296 -57 314 -55 0 FreeSans 56 0 0 -56 V2
flabel metal1 465 -69 481 -67 0 FreeSans 56 0 0 -56 V3
flabel metal1 298 -152 314 -150 0 FreeSans 56 0 0 -56 V4
flabel metal1 -45 547 -42 564 0 FreeSans 40 90 0 56 VOUT1
flabel metal1 651 547 653 564 0 FreeSans 40 270 0 56 VOUT2
<< end >>
